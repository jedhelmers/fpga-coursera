/*
  74LS161a replacement
  4-bit binary counter
  for Coursera course: Hardware Description Languages

  D:        Parallel Input
  CLK:      Clock
  CLR_n:    Asynchronous Reset (LOW)
  LOAD_n:   Enable Parallel Input (LOW)
  ENP:      Count Enable Parallel
  ENT:      Count Enable Trickle
  Q:        Parallel Output
  RCO:      Ripple Carry Output (Terminal Count)

*/
module LS161a(
    input [3:0] D,
    input CLK,
    input CLR_n,
    input LOAD_n,
    input ENP,
    input ENT,
    output RCO,
    output [3:0]Q
);
  reg [4:0] CNT;

  assign Q = CNT[3:0];

  assign RCO = CNT[4];

  always @(posedge CLK or negedge LOAD_n) begin
    if (!LOAD_n) begin
      $display("!LOAD_n: D %d Q %d", D, Q);
      CNT = D;
    end
  end

  always @(posedge CLK or posedge CLR_n) begin
    if (!CLR_n) begin
      CNT <= 0;
    end
    else begin
      if (ENP) begin
        CNT = CNT + 1;
        $display("%b", CNT);
      end
      if(CNT > 5'b10000) begin
        CNT <= 0;
      end
    end
  end
endmodule